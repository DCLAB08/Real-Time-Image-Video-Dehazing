
module VGA_pll (
	clk_clk,
	clk_120m_clk,
	clk_100m_clk,
	clk_75m_clk,
	clk_800k_clk,
	reset_reset_n);	

	input		clk_clk;
	output		clk_120m_clk;
	output		clk_100m_clk;
	output		clk_75m_clk;
	output		clk_800k_clk;
	input		reset_reset_n;
endmodule
